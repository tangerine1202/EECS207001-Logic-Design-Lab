`timescale 1ns/1ps

module Carry_Look_Ahead_Adder_t;

endmodule
