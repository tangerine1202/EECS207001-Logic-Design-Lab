`timescale 1ns/1ps

module LFSR (clk, rst_n, out);
input clk, rst_n;
output out;

endmodule
